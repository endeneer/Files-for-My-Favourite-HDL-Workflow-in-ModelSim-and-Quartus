module myxorgate
    (
    input  i_A,
    input  i_B,
    output o_C
    );

    assign o_C = i_A ^ i_B;
endmodule
